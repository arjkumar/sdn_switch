library verilog;
use verilog.vl_types.all;
entity header_hash_tester is
end header_hash_tester;
